-- TI Proprietary Information - Internal Data.  Copyright (c) 2011, Texas Instruments Incorporated.  All rights reserved.
library IEEE; use IEEE.Std_Logic_1164.all; use IEEE.Std_Logic_arith.all; use IEEE.Std_Logic_unsigned.all; library work; use work.dtsa_cj_pkg.all; entity dtsa_tclk_ctrl is port(reset_n:in std_logic; reset_n_fe:in std_logic; master_clk:in std_logic; wr_clr_det:in std_logic; 
ctr_limit:in std_logic_vector(5 downto 0); tck_cfg_mode:in std_logic_vector(K29 downto K30); clk_1500:in std_logic; jscan_fmt:in std_logic; csm_to_std:in std_logic; ts_rtck_pin:in std_logic; ctlr_tck_pin:in std_logic; tck_en:in std_logic; tap_adv:in std_logic; csm_std_mode:in std_logic; csm_run:in std_logic; 
clr_clk_fail:in std_logic; clk_fail:out std_logic; clk_det:out std_logic; clk_tst:out std_logic; ctlr_rtck:out std_logic; tck2tgt:out std_logic; itck:out std_logic ); end dtsa_tclk_ctrl; architecture RTL of dtsa_tclk_ctrl is CONSTANT ITCK_BIT:integer:=3; 
CONSTANT TCK_BIT:integer:=2; CONSTANT RTCK_BIT:integer:=1; CONSTANT CLK_LO_ST:std_logic_vector(3 downto 0):="0000"; CONSTANT STD_HI_ST:std_logic_vector(3 downto 0):="1101"; CONSTANT RTCK_HI_ST:std_logic_vector(3 downto 0):="1111"; CONSTANT RTCK_LO_ST:std_logic_vector(3 downto 0):="0010"; CONSTANT ADV_HI_ST:std_logic_vector(3 downto 0):="1100"; CONSTANT ADV_LO_ST:std_logic_vector(3 downto 0):="0001"; CONSTANT ESC_LO_ST:std_logic_vector(3 downto 0):="0100"; CONSTANT ADV_END_ST:std_logic_vector(3 downto 0):="0011"; CONSTANT CP_END_ST:std_logic_vector(3 downto 0):="1001"; 
signal tsm_pres_st:std_logic_vector(3 downto 0); signal tsm_next_st:std_logic_vector(3 downto 0); signal clr_clk_fail_r:std_logic; signal clk_det_in:std_logic; signal clk_det_hi:std_logic; signal clk_det_lo:std_logic; signal clk_fail_in:std_logic; signal clk_fail_r:std_logic; signal clk_timeout:std_logic; signal csm_run_flg:std_logic; signal csm_run_dly:std_logic; 
signal csm_start:std_logic; signal csm_start_mode:std_logic; signal ctlr_tck_sync:std_logic; signal ctr_eq_1:std_logic; signal ctr_eq_0_q:std_logic; signal ctr_lim_eq_0:std_logic; signal free_run_mode:std_logic; signal level_ctr:std_logic_vector(1 downto 0); signal level_ctr_is_3:std_logic; signal limit_eq_0:std_logic; signal mismatch:std_logic; 
signal mismatch_ctr:std_logic_vector(1 downto 0); signal mm_ctr_is_3:std_logic; signal rtck_re:std_logic; signal rtck_sync:std_logic; signal rtck_sync2:std_logic; signal same_level:std_logic; signal std_2_adv:std_logic; signal tck_ctr:std_logic_vector(5 downto 0); signal tck_re:std_logic; signal tck_sync:std_logic; signal tck_sync2:std_logic; 
signal tck_sync_mode:std_logic; signal ts_rtck_sync:std_logic; signal tck_sync_lo:std_logic; signal tck_sync_hi:std_logic; begin tck_sync_mode<='1'when tck_cfg_mode=K33 else'0'; free_run_mode<='1'when tck_cfg_mode=K32 else'0'; I33:process(reset_n_fe,master_clk) begin if(reset_n_fe='0')then ctlr_tck_sync<='0'; 
elsif(master_clk'event and master_clk='0')then ctlr_tck_sync<=ctlr_tck_pin; end if; end process I33; I34:process(reset_n,master_clk) begin if(reset_n='0')then tck_sync<='0'; tck_sync2<='0'; elsif(master_clk'event and master_clk='1')then tck_sync<=ctlr_tck_sync; 
tck_sync2<=tck_sync; end if; end process I34; I35:process(reset_n,master_clk) begin if(reset_n='0')then tck_sync_lo<='0'; tck_sync_hi<='0'; elsif(master_clk'event and master_clk='1')then tck_sync_lo<=not ctlr_tck_sync OR free_run_mode; tck_sync_hi<=ctlr_tck_sync OR free_run_mode; 
end if; end process I35; tck_re<=tck_sync AND not tck_sync2; I36:process(reset_n_fe,master_clk) begin if(reset_n_fe='0')then ts_rtck_sync<='0'; elsif(master_clk'event and master_clk='0')then ts_rtck_sync<=ts_rtck_pin; end if; end process I36; 
I37:process(reset_n,master_clk) begin if(reset_n='0')then rtck_sync<='0'; elsif(master_clk'event and master_clk='1')then rtck_sync<=ts_rtck_sync; end if; end process I37; I38:process(reset_n,master_clk) begin if(reset_n='0')then 
rtck_sync2<='0'; elsif(master_clk'event and master_clk='1')then rtck_sync2<=tsm_pres_st(RTCK_BIT); end if; end process I38; rtck_re<=tsm_pres_st(RTCK_BIT)AND not rtck_sync2; limit_eq_0<='1'when ctr_limit="000000"else'0'; process(reset_n,master_clk) begin if(reset_n='0')then ctr_lim_eq_0<='0'; 
elsif(master_clk'event and master_clk='1')then ctr_lim_eq_0<=limit_eq_0; end if; end process; I39:process(reset_n,master_clk) begin if(reset_n='0')then tck_ctr<="000000"; elsif(master_clk'event and master_clk='1')then if(ctr_eq_0_q='1')then tck_ctr<=ctr_limit; 
else tck_ctr<=tck_ctr-"000001"; end if; end if; end process I39; ctr_eq_1<='1'when tck_ctr="000001"else'0'; I40:process(reset_n,master_clk) begin if(reset_n='0')then ctr_eq_0_q<='0'; elsif(master_clk'event and master_clk='1')then 
ctr_eq_0_q<=ctr_eq_1 OR ctr_lim_eq_0; end if; end process I40; I41:process(master_clk,reset_n) begin if(reset_n='0')then tsm_pres_st<=CLK_LO_ST; elsif(master_clk'event AND master_clk='1')then if(ctr_eq_0_q='1')then tsm_pres_st<=tsm_next_st; end if; 
end if; end process I41; tck2tgt<=tsm_pres_st(TCK_BIT); ctlr_rtck<=tsm_pres_st(RTCK_BIT); itck<=tsm_pres_st(ITCK_BIT); I42:process(master_clk,reset_n) begin if(reset_n='0')then clk_tst<='0'; elsif(master_clk'event AND master_clk='1')then clk_tst<=ctr_eq_1 OR ctr_lim_eq_0; 
end if; end process I42; process(master_clk,reset_n) begin if(reset_n='0')then csm_run_dly<='0'; elsif(master_clk'event AND master_clk='1')then csm_run_dly<=csm_run; end if; end process; csm_start<=csm_run AND not csm_run_dly; 
process(master_clk,reset_n) begin if(reset_n='0')then csm_start_mode<='0'; elsif(master_clk'event AND master_clk='1')then if(csm_start='1')then csm_start_mode<=csm_std_mode; end if; end if; end process; std_2_adv<=csm_start_mode AND not jscan_fmt; 
process(master_clk,reset_n) begin if(reset_n='0')then csm_run_flg<='0'; elsif(master_clk'event AND master_clk='1')then if(tsm_pres_st=CLK_LO_ST)then csm_run_flg<='0'; else csm_run_flg<=(csm_run OR csm_run_flg)AND std_2_adv; end if; end if; 
end process; process(tsm_pres_st,tck_sync_lo,tck_sync_hi,csm_std_mode,rtck_sync, tck_sync_mode,csm_run,tap_adv,tck_en,csm_to_std,csm_run_flg) begin CASE tsm_pres_st IS WHEN CLK_LO_ST=> if(tck_sync_hi AND(csm_run OR not csm_std_mode))='1'then tsm_next_st<=ADV_HI_ST; elsif(tck_sync_hi AND csm_std_mode)='1'then tsm_next_st<=STD_HI_ST; else 
tsm_next_st<=CLK_LO_ST; end if; WHEN STD_HI_ST=> if(rtck_sync='1')OR(tck_sync_mode='1')then tsm_next_st<=RTCK_HI_ST; else tsm_next_st<=STD_HI_ST; end if; WHEN RTCK_HI_ST=> if(tck_sync_lo='1')then tsm_next_st<=RTCK_LO_ST; 
else tsm_next_st<=RTCK_HI_ST; end if; WHEN RTCK_LO_ST=> if(rtck_sync='0')OR(tck_sync_mode='1')then tsm_next_st<=CLK_LO_ST; else tsm_next_st<=RTCK_LO_ST; end if; WHEN ADV_HI_ST=> if(tck_en='0')OR(csm_to_std='1')then 
tsm_next_st<=ESC_LO_ST; else tsm_next_st<=ADV_LO_ST; end if; WHEN ADV_LO_ST=> if(csm_run='0'AND tap_adv='1')then if(csm_run_flg='1')then tsm_next_st<=CP_END_ST; else tsm_next_st<=ADV_END_ST; end if; 
else tsm_next_st<=ADV_HI_ST; end if; WHEN ESC_LO_ST=> tsm_next_st<=ADV_HI_ST; WHEN ADV_END_ST=> if(tck_sync_lo='1')then tsm_next_st<=CLK_LO_ST; else tsm_next_st<=ADV_END_ST; end if; 
WHEN CP_END_ST=> tsm_next_st<=RTCK_HI_ST; WHEN others=> tsm_next_st<=CLK_LO_ST; END CASE; end process; I43:process(reset_n,master_clk) begin if(reset_n='0')then clk_det_in<='0'; elsif(master_clk'event and master_clk='1')then 
clk_det_in<=ts_rtck_pin; end if; end process I43; I44:process(reset_n,master_clk) begin if(reset_n='0')then clk_det_hi<='0'; elsif(master_clk'event and master_clk='1')then clk_det_hi<=(clk_det_in OR clk_det_hi)AND not wr_clr_det; end if; end process I44; 
I45:process(reset_n,master_clk) begin if(reset_n='0')then clk_det_lo<='0'; elsif(master_clk'event and master_clk='1')then clk_det_lo<=(not clk_det_in OR clk_det_lo)AND not wr_clr_det; end if; end process I45; I46:process(reset_n,master_clk) begin if(reset_n='0')then 
clk_det<='0'; elsif(master_clk'event and master_clk='1')then clk_det<=clk_det_lo AND clk_det_hi AND not wr_clr_det; end if; end process I46; process(master_clk,reset_n) begin if(reset_n='0')then clr_clk_fail_r<='1'; elsif(master_clk'event AND master_clk='1')then clr_clk_fail_r<=(clr_clk_fail OR clr_clk_fail_r)AND not rtck_re; 
end if; end process; process(master_clk,reset_n) begin if(reset_n='0')then mismatch_ctr<="00"; elsif(master_clk'event AND master_clk='1')then if(clr_clk_fail_r='1')then mismatch_ctr<="00"; elsif(tck_re='1')AND(rtck_re='0')then mismatch_ctr<=mismatch_ctr+"01"; 
elsif(tck_re='0')AND(rtck_re='1')then mismatch_ctr<=mismatch_ctr-"01"; end if; end if; end process; mm_ctr_is_3<='1'when mismatch_ctr="11"else'0'; process(master_clk,reset_n) begin if(reset_n='0')then mismatch<='0'; elsif(master_clk'event AND master_clk='1')then 
mismatch<=mm_ctr_is_3; end if; end process; same_level<=not(tck_sync XOR tsm_pres_st(RTCK_BIT)); process(master_clk,reset_n) begin if(reset_n='0')then level_ctr<="00"; elsif(master_clk'event AND master_clk='1')then if(clr_clk_fail='1')or(same_level='1')then level_ctr<="00"; 
elsif(clk_1500='1')then level_ctr<=level_ctr+"01"; end if; end if; end process; level_ctr_is_3<='1'when level_ctr="11"else'0'; process(master_clk,reset_n) begin if(reset_n='0')then clk_timeout<='0'; elsif(master_clk'event AND master_clk='1')then 
clk_timeout<=level_ctr_is_3; end if; end process; clk_fail_in<=(clk_fail_r OR clk_timeout OR mismatch)AND not clr_clk_fail; process(master_clk,reset_n) begin if(reset_n='0')then clk_fail_r<='0'; elsif(master_clk'event AND master_clk='1')then clk_fail_r<=clk_fail_in; end if; 
end process; clk_fail<=clk_fail_r; end RTL; 