-- TI Proprietary Information - Internal Data.  Copyright (c) 2011, Texas Instruments Incorporated.  All rights reserved.
library ieee; use ieee.std_logic_1164.all; package dtsa_cj_pkg is constant K0:std_logic_vector(7 downto 4):="0001"; constant K1:std_logic_vector(7 downto 4):="0010"; constant K2:std_logic_vector(7 downto 4):="0011"; constant K3:std_logic_vector(7 downto 4):="0100"; constant K4:std_logic_vector(7 downto 4):="0101"; constant K5:std_logic_vector(3 downto 0):="0001"; constant K6:std_logic_vector(7 downto 0):=X"5A"; constant K7:std_logic_vector(31 downto 0):=X"00000000"; 
constant K8:integer:=7; constant K9:std_logic_vector(7 downto 0):="00000000"; constant K10:std_logic_vector(7 downto 0):="00000001"; constant K11:std_logic_vector(7 downto 0):="00000010"; constant K12:std_logic_vector(7 downto 0):="00000011"; constant K13:std_logic_vector(7 downto 0):="00000100"; constant K14:std_logic_vector(7 downto 0):="00000101"; constant K15:std_logic_vector(7 downto 0):="00000110"; constant K16:std_logic_vector(7 downto 0):="00000111"; constant K17:std_logic_vector(7 downto 0):="00001000"; constant K18:std_logic_vector(7 downto 0):="00000001"; 
constant K19:integer:=7; constant K20:integer:=6; constant K21:integer:=5; constant K22:integer:=4; constant K23:integer:=128; constant K24:integer:=64; constant K25:integer:=32; constant K26:integer:=16; constant K27:integer:=5; constant K28:integer:=0; constant K29:integer:=2; 
constant K30:integer:=0; constant K31:std_logic_vector(2 downto 0):="101"; constant K32:std_logic_vector(2 downto 0):="100"; constant K33:std_logic_vector(2 downto 0):="000"; constant K34:integer:=5; constant K35:integer:=4; constant K36:integer:=0; constant K37:integer:=7; constant K38:integer:=6; constant K39:integer:=5; constant K40:integer:=4; 
constant K41:integer:=3; constant K42:integer:=2; constant K43:integer:=1; constant K44:integer:=0; constant K45:integer:=1; constant K46:integer:=0; constant K47:integer:=2; constant K48:integer:=1; constant K49:integer:=7; constant K50:integer:=6; constant K51:integer:=5; 
constant K52:integer:=4; constant K53:integer:=3; constant K54:integer:=1; constant K55:integer:=0; constant K56:integer:=7; constant K57:integer:=5; constant K58:integer:=4; constant K59:integer:=3; constant K60:integer:=2; constant K61:integer:=1; constant K62:integer:=0; 
constant K63:integer:=9; constant K64:std_logic_vector(9 downto 0):="0010000001"; constant K65:std_logic_vector(9 downto 0):="0010000010"; constant K66:std_logic_vector(9 downto 0):="0010000100"; constant K67:std_logic_vector(9 downto 0):="0010001000"; constant K68:std_logic_vector(9 downto 0):="0010010000"; constant K69:std_logic_vector(9 downto 0):="0010100000"; constant K70:std_logic_vector(9 downto 0):="0011000000"; constant K71:std_logic_vector(9 downto 0):="0000000001"; constant K72:std_logic_vector(9 downto 0):="0000000010"; constant K73:std_logic_vector(9 downto 0):="0000000100"; 
constant K74:std_logic_vector(9 downto 0):="0000001000"; constant K75:std_logic_vector(9 downto 0):="0000010000"; constant K76:std_logic_vector(9 downto 0):="0000100000"; constant K77:std_logic_vector(9 downto 0):="0001000000"; constant K78:std_logic_vector(9 downto 0):="0100000000"; constant K79:std_logic_vector(9 downto 0):="1000000000"; constant K80:integer:=0; constant K81:integer:=1; constant K82:integer:=2; constant K83:integer:=3; constant K84:integer:=4; 
constant K85:integer:=5; constant K86:integer:=6; constant K87:integer:=7; constant K88:integer:=8; constant K89:integer:=9; constant K90:std_logic_vector(3 downto 0):="0000"; constant K91:std_logic_vector(3 downto 0):="1000"; constant K92:std_logic_vector(3 downto 0):="0001"; constant K93:std_logic_vector(3 downto 0):="0010"; constant K94:std_logic_vector(3 downto 0):="0011"; constant K95:std_logic_vector(3 downto 0):="0100"; 
constant K96:std_logic_vector(3 downto 0):="0101"; constant K97:std_logic_vector(3 downto 0):="0110"; constant K98:std_logic_vector(3 downto 0):="0111"; constant K99:std_logic_vector(3 downto 0):="1001"; constant K100:std_logic_vector(3 downto 0):="1010"; constant K101:std_logic_vector(3 downto 0):="1011"; constant K102:std_logic_vector(3 downto 0):="1100"; constant K103:std_logic_vector(3 downto 0):="1101"; constant K104:std_logic_vector(3 downto 0):="1110"; constant K105:std_logic_vector(3 downto 0):="1111"; constant K106:integer:=4; 
constant K107:integer:=4; constant K108:integer:=9; constant K109:std_logic_vector(4 downto 0):="00000"; constant K110:std_logic_vector(4 downto 0):="00001"; constant K111:std_logic_vector(4 downto 0):="00010"; constant K112:std_logic_vector(4 downto 0):="00011"; constant K113:std_logic_vector(4 downto 0):="00100"; constant K114:std_logic_vector(4 downto 0):="00101"; constant K115:std_logic_vector(4 downto 0):="00110"; constant K116:std_logic_vector(4 downto 0):="00111"; constant K117:std_logic_vector(4 downto 0):="01000"; 
constant K118:std_logic_vector(4 downto 0):="01001"; constant K119:std_logic_vector(4 downto 0):="01010"; constant K120:std_logic_vector(4 downto 0):="01011"; constant K121:std_logic_vector(4 downto 0):="00001"; constant K122:std_logic_vector(4 downto 2):="010"; constant K123:std_logic_vector(4 downto 2):="011"; constant K124:std_logic_vector(4 downto 2):="101"; constant K125:std_logic_vector(4 downto 2):="110"; constant K126:std_logic_vector(3 downto 0):="1001"; constant K127:std_logic_vector(4 downto 0):="00111"; constant K128:std_logic_vector(2 downto 0):="000"; 
constant K129:integer:=4; constant K130:std_logic_vector(4 downto 0):="00000"; constant K131:std_logic_vector(4 downto 0):="00001"; constant K132:std_logic_vector(4 downto 0):="00010"; constant K133:std_logic_vector(4 downto 0):="00011"; constant K134:std_logic_vector(4 downto 0):="00100"; constant K135:std_logic_vector(4 downto 0):="00101"; constant K136:std_logic_vector(4 downto 0):="00110"; constant K137:std_logic_vector(4 downto 0):="00111"; constant K138:std_logic_vector(4 downto 0):="01000"; constant K139:std_logic_vector(4 downto 0):="01001"; 
constant K140:std_logic_vector(4 downto 0):="01010"; constant K141:std_logic_vector(4 downto 0):="01011"; constant K142:std_logic_vector(4 downto 0):="01100"; constant K143:std_logic_vector(4 downto 0):="01101"; constant K144:std_logic_vector(4 downto 0):="01110"; constant K145:std_logic_vector(4 downto 0):="01111"; constant K146:std_logic_vector(4 downto 0):="10000"; constant K147:integer:=0; constant K148:integer:=1; constant K149:integer:=2; constant K150:integer:=3; 
constant K151:integer:=4; constant K152:integer:=5; constant K153:integer:=6; constant K154:integer:=7; constant K155:integer:=8; constant K156:integer:=9; constant K157:integer:=9; constant K158:integer:=5; constant K159:std_logic_vector(5 downto 0):="000001"; constant K160:std_logic_vector(5 downto 0):="000010"; constant K161:std_logic_vector(5 downto 0):="000100"; 
constant K162:std_logic_vector(5 downto 0):="001000"; constant K163:std_logic_vector(5 downto 0):="010000"; constant K164:std_logic_vector(5 downto 0):="100000"; constant K165:integer:=0; constant K166:integer:=1; constant K167:integer:=2; constant K168:integer:=3; constant K169:integer:=4; constant K170:integer:=5; end package dtsa_cj_pkg; 